`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/10/27 09:37:19
// Design Name: 
// Module Name: rotword_subword_rcon_with_smaller_area
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rotword_subword_rcon_with_smaller_area(
    input   [31:0]      input_data,
    input   [1:0]       key_width,                          //2'b00 means 128bit ,2'b01 means 192bit, 2'b10 means 256bit
    
  /*  
    input   [2:0]       key_expand_cycle_number,            //cycle_number record which cycle in one round,when cycle_number = 3'b0,need rotword+subword+rcon;when cycle_number = 3'd4,need subword
  */  
    
    input   [3:0]       key_expand_round_number,            //round number record which round
    input   [1:0]       control_signal,                     //this signal is generated by key expansion module
                                                            //2'b00 means default, 2'b01 means sbox with rcon and shiftrow, 2'b10 means only sbox
    output  [31:0]      output_data
    );
    
    wire    [31:0]      w0,w1,w2,w3,w4;
    wire    [7:0]       rcon;
    
    assign   w0 =   input_data;
    assign   w1 =   w3;
    assign   w4 =   {w3[23:16],w3[15:08],w3[07:00],w3[31:24]};      //rotword
    assign   w2 =   {w4[31:24]^rcon,w4[23:0]};
    
    assign   output_data    =   (control_signal == 2'b01) ? w2 : (control_signal == 2'b10) ? w1 : w0;
    
    sbox_in_GF16_with_only_affine       u0_sbox_in_GF16_with_only_affine(
    .input_of_inv_and_affine_in_GF16    (input_data[31:24]),
    .output_of_inv_and_affine_in_GF16   (w3[31:24])
    );
    
    sbox_in_GF16_with_only_affine       u1_sbox_in_GF16_with_only_affine(
    .input_of_inv_and_affine_in_GF16    (input_data[23:16]),
    .output_of_inv_and_affine_in_GF16   (w3[23:16])
    );
    
    sbox_in_GF16_with_only_affine       u2_sbox_in_GF16_with_only_affine(
    .input_of_inv_and_affine_in_GF16    (input_data[15:08]),
    .output_of_inv_and_affine_in_GF16   (w3[15:08])
    );
    
    sbox_in_GF16_with_only_affine       u3_sbox_in_GF16_with_only_affine(
    .input_of_inv_and_affine_in_GF16    (input_data[07:00]),
    .output_of_inv_and_affine_in_GF16   (w3[07:00])
    );
        
    rcon                    u_rcon(
    .key_expand_round_number    (key_expand_round_number),
    .rcon                       (rcon)
    );
endmodule
